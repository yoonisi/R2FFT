�� 
 m o d u l e   t w i d d l e F a c t o r R o m B r i d g e  
     # (  
         p a r a m e t e r   F F T _ N   =   1 0 ,  
         p a r a m e t e r   F F T _ D W   =   1 6  
         )  
     (  
       i n p u t   w i r e                                       c l k ,  
       i n p u t   w i r e                                       r s t ,  
       i n p u t   w i r e                                       t a c t _ r o m ,  
       i n p u t   w i r e   [ F F T _ N - 1 - 1 : 0 ]           t a _ r o m ,  
  
       i n p u t   w i r e                                       e v e n O d d ,  
       i n p u t   w i r e                                       i f f t ,  
        
       o u t p u t   r e g   s i g n e d   [ F F T _ D W : 0 ]   t d r _ r o m _ r e a l ,  
       o u t p u t   r e g   s i g n e d   [ F F T _ D W : 0 ]   t d r _ r o m _ i m a g ,  
  
       / /   t w i d d l e   f a c t o r   r o m   i n t e r f a c e  
       o u t p u t   w i r e                                     t w a c t ,  
       o u t p u t   w i r e   [ F F T _ N - 1 - 2 : 0 ]         t w a ,  
       i n p u t   w i r e   [ F F T _ D W - 1 : 0 ]         t w d r _ c o s  
       ) ;  
  
  
       / /   p i p e l i n e   s t a g e   1  
       r e g                                             t a c t _ 1 ;  
       r e g                                             t a _ m s b _ 1 ;  
       w i r e   [ F F T _ N - 1 - 2 : 0 ]               c o s A d d r   =   t a _ r o m [ F F T _ N - 1 - 2 : 0 ] ;  
       r e g                                             e v e n O d d _ 1 ;  
       / /   p i p e l i n e   s t a g e   2  
       r e g   [ F F T _ N - 1 - 2 : 0 ]   	         s i n A d d r ;  
       r e g                                             t a c t _ 2 ;  
       r e g                                             t a _ m s b _ 2 ;  
       r e g                                             e v e n O d d _ 2 ;  
  
       / /   p i p e l i n e   s t a g e   3  
       r e g                                             t a _ m s b _ 3 ;  
  
       a l w a y s   @   (   p o s e d g e   c l k   )   b e g i n  
             i f   (   r s t   )   b e g i n  
                   t a c t _ 1   < =   0 ;  
                   t a _ m s b _ 1   < =   0 ;  
                   s i n A d d r   < =   0 ;  
                   e v e n O d d _ 1   < =   0 ;  
                    
                   t a c t _ 2   < =   0 ;  
                   t a _ m s b _ 2   < =   0 ;  
                   e v e n O d d _ 2   < =   0 ;  
  
                   t a _ m s b _ 3   < =   0 ;  
             e n d   e l s e   b e g i n  
                    
                   t a c t _ 1   < =   t a c t _ r o m ;  
                   t a _ m s b _ 1   < =   t a _ r o m [ F F T _ N - 1 - 1 ] ;  
                   s i n A d d r   < =   { 1 ' b 1 , { ( F F T _ N - 1 - 1 ) { 1 ' b 0 } } }   -   t a _ r o m [ F F T _ N - 1 - 2 : 0 ] ;  
                   e v e n O d d _ 1   < =   e v e n O d d ;  
                    
                   t a c t _ 2   < =   t a c t _ 1 ;  
                   t a _ m s b _ 2   < =   t a _ m s b _ 1 ;  
                   e v e n O d d _ 2   < =   e v e n O d d _ 1 ;  
  
                   t a _ m s b _ 3   < =   t a _ m s b _ 2 ;  
             e n d  
       e n d   / /   a l w a y s   @   (   p o s e d g e   c l k   )  
  
       w i r e   c o s R o m A d d r P h a s e   =   t a c t _ r o m   & &   ( e v e n O d d   = =   1 ' b 0 ) ;  
       w i r e   c o s R o m D a t a P h a s e   =   t a c t _ 1       & &   ( e v e n O d d _ 1   = =   1 ' b 0 ) ;  
       w i r e   s i n R o m A d d r P h a s e   =   c o s R o m D a t a P h a s e ;  
       w i r e   s i n R o m D a t a P h a s e   =   t a c t _ 2       & &   ( e v e n O d d _ 2   = =   1 ' b 0 ) ;  
  
       a s s i g n   t w a c t   =   c o s R o m A d d r P h a s e   | |   s i n R o m A d d r P h a s e ;  
       a s s i g n   t w a       =   s i n R o m A d d r P h a s e   ?   s i n A d d r   :   c o s A d d r ;  
  
       r e g   	 s i n 0 ;  
       a l w a y s   @   (   p o s e d g e   c l k   )   b e g i n  
             s i n 0   < =   (   s i n A d d r   = =   0   )   ?   1 ' b 1   :   1 ' b 0 ;  
       e n d  
        
       w i r e   s i g n e d   [ F F T _ D W : 0 ]   c o s R e a d D a t a   =   { 1 ' b 0 ,   t w d r _ c o s } ;  
       w i r e   s i g n e d   [ F F T _ D W : 0 ]   s i n R e a d D a t a   =   s i n 0   ?   0   :   { 1 ' b 0 ,   t w d r _ c o s } ;  
  
       r e g   s i g n e d   [ F F T _ D W : 0 ]     c o s R e a d D a t a _ 1 ;  
       r e g   s i g n e d   [ F F T _ D W : 0 ]     c o s R e a d D a t a _ 2 ;  
       a l w a y s   @   (   p o s e d g e   c l k   )   b e g i n  
             i f   (   c o s R o m D a t a P h a s e   )   b e g i n  
                   c o s R e a d D a t a _ 1   < =   c o s R e a d D a t a ;  
             e n d  
             c o s R e a d D a t a _ 2   < =   c o s R e a d D a t a _ 1 ;  
       e n d  
  
       r e g   s i g n e d   [ F F T _ D W : 0 ]   s i n R e a d D a t a _ 2 ;  
       a l w a y s   @   (   p o s e d g e   c l k   )   b e g i n  
             i f   (   s i n R o m D a t a P h a s e   )   b e g i n  
                   s i n R e a d D a t a _ 2   < =   s i n R e a d D a t a ;  
             e n d  
       e n d  
  
       a l w a y s _ c o m b   b e g i n  
             i f   (   t a _ m s b _ 3   = =   1 ' b 0   )   b e g i n  
                   t d r _ r o m _ r e a l   =   c o s R e a d D a t a _ 2 ;  
                   t d r _ r o m _ i m a g   =   i f f t   ?   s i n R e a d D a t a _ 2   :   - s i n R e a d D a t a _ 2 ;  
             e n d   e l s e   b e g i n  
                   t d r _ r o m _ r e a l   =   - s i n R e a d D a t a _ 2 ;  
                   t d r _ r o m _ i m a g   =   i f f t   ?   c o s R e a d D a t a _ 2   :   - c o s R e a d D a t a _ 2 ;  
             e n d  
       e n d  
        
 e n d m o d u l e   / /   t w i d d l e F a c t o r R o m  
  
 